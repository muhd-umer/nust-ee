** Profile: "SCHEMATIC1-A"  [ D:\NUST\SEMESTER 4\ELECTRONIC DEVICES AND CIRCUITS\LABS\Lab 10\lab10-SCHEMATIC1-A.sim ] 

** Creating circuit file "lab10-SCHEMATIC1-A.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10m 0 0.00001 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\lab10-SCHEMATIC1.net" 


.END
