** Profile: "SCHEMATIC1-Lab"  [ F:\NUST\Semester 1\Linear Circuit Analysis\Labs\PSpice\apl3-SCHEMATIC1-Lab.sim ] 

** Creating circuit file "apl3-SCHEMATIC1-Lab.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\apl3-SCHEMATIC1.net" 


.END
