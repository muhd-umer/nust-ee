** Profile: "SCHEMATIC1-asd"  [ F:\NUST\Semester 1\Linear Circuit Analysis\Labs\PSpice\lab11and12-schematic1-asd.sim ] 

** Creating circuit file "lab11and12-schematic1-asd.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 40ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\lab11and12-SCHEMATIC1.net" 


.END
