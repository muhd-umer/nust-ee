** Profile: "SCHEMATIC1-f"  [ F:\NUST\Semester 1\Linear Circuit Analysis\Labs\PSpice\op-SCHEMATIC1-f.sim ] 

** Creating circuit file "op-SCHEMATIC1-f.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\op-SCHEMATIC1.net" 


.END
