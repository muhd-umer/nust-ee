** Profile: "SCHEMATIC1-A"  [ F:\NUST\Semester 2\Electric Network Analysis\PSpice\lab 4-SCHEMATIC1-A.sim ] 

** Creating circuit file "lab 4-SCHEMATIC1-A.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 50m 0 0.005m 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\lab 4-SCHEMATIC1.net" 


.END
