** Profile: "SCHEMATIC1-a"  [ F:\NUST\Semester 1\Linear Circuit Analysis\Labs\PSpice\asddfg-SCHEMATIC1-a.sim ] 

** Creating circuit file "asddfg-SCHEMATIC1-a.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\asddfg-SCHEMATIC1.net" 


.END
