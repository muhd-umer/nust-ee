** Profile: "SCHEMATIC1-sasd"  [ F:\NUST\Semester 1\Linear Circuit Analysis\Labs\PSpice\quiz1-SCHEMATIC1-sasd.sim ] 

** Creating circuit file "quiz1-SCHEMATIC1-sasd.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\quiz1-SCHEMATIC1.net" 


.END
