** Profile: "SCHEMATIC1-s"  [ F:\NUST\Semester 1\Linear Circuit Analysis\Labs\PSpice\quiz-SCHEMATIC1-s.sim ] 

** Creating circuit file "quiz-SCHEMATIC1-s.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\quiz-SCHEMATIC1.net" 


.END
