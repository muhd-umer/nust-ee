** Profile: "SCHEMATIC1-ad"  [ F:\NUST\Semester 1\Linear Circuit Analysis\Labs\PSpice\exam-SCHEMATIC1-ad.sim ] 

** Creating circuit file "exam-SCHEMATIC1-ad.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\exam-SCHEMATIC1.net" 


.END
