** Profile: "SCHEMATIC1-fdg"  [ F:\NUST\Semester 1\Linear Circuit Analysis\Labs\PSpice\yui-SCHEMATIC1-fdg.sim ] 

** Creating circuit file "yui-SCHEMATIC1-fdg.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\yui-SCHEMATIC1.net" 


.END
