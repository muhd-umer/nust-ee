** Profile: "SCHEMATIC1-a"  [ D:\NUST\SEMESTER 4\ELECTRONIC DEVICES AND CIRCUITS\LABS\Lab 4\lab4-schematic1-a.sim ] 

** Creating circuit file "lab4-schematic1-a.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 50m 0 2u 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\lab4-SCHEMATIC1.net" 


.END
