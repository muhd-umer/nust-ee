** Profile: "SCHEMATIC1-ASD"  [ F:\NUST\Semester 1\Linear Circuit Analysis\Labs\PSpice\lab1112-SCHEMATIC1-ASD.sim ] 

** Creating circuit file "lab1112-SCHEMATIC1-ASD.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 80m 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\lab1112-SCHEMATIC1.net" 


.END
