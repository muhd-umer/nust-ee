** Profile: "SCHEMATIC1-sa"  [ D:\NUST\SEMESTER 4\ELECTRONIC DEVICES AND CIRCUITS\LABS\Lab 4\lab4-SCHEMATIC1-sa.sim ] 

** Creating circuit file "lab4-SCHEMATIC1-sa.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 50ms 0 2u 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\lab4-SCHEMATIC1.net" 


.END
