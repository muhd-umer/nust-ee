** Profile: "SCHEMATIC1-b"  [ D:\NUST\SEMESTER 4\ELECTRONIC DEVICES AND CIRCUITS\LABS\Lab 5\main-SCHEMATIC1-b.sim ] 

** Creating circuit file "main-SCHEMATIC1-b.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V3 0 10 0.2 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\main-SCHEMATIC1.net" 


.END
