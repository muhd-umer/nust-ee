** Profile: "SCHEMATIC3-task3"  [ D:\NUST\Semester 4\Electronic Devices and Circuits\Labs\Lab 1\lab1-schematic3-task3.sim ] 

** Creating circuit file "lab1-schematic3-task3.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\lab1-SCHEMATIC3.net" 


.END
