** Profile: "SCHEMATIC1-sd"  [ F:\NUST\Semester 1\Linear Circuit Analysis\Labs\PSpice\asd-SCHEMATIC1-sd.sim ] 

** Creating circuit file "asd-SCHEMATIC1-sd.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\asd-SCHEMATIC1.net" 


.END
