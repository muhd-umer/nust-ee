** Profile: "SCHEMATIC1-A"  [ F:\NUST\Semester 1\Linear Circuit Analysis\Labs\PSpice\lab6-SCHEMATIC1-A.sim ] 

** Creating circuit file "lab6-SCHEMATIC1-A.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\lab6-SCHEMATIC1.net" 


.END
