** Profile: "SCHEMATIC1-a"  [ D:\NUST\Semester 1\Linear Circuit Analysis\Labs\PSpice\a-schematic1-a.sim ] 

** Creating circuit file "a-schematic1-a.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\a-SCHEMATIC1.net" 


.END
