** Profile: "SCHEMATIC2-task2"  [ D:\NUST\Semester 4\Electronic Devices and Circuits\Labs\Lab 1\lab1-SCHEMATIC2-task2.sim ] 

** Creating circuit file "lab1-SCHEMATIC2-task2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V1 0 20 0.1 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\lab1-SCHEMATIC2.net" 


.END
