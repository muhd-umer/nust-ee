** Profile: "SCHEMATIC1-Sim"  [ D:\NUST\SEMESTER 4\ELECTRONIC DEVICES AND CIRCUITS\LABS\Lab 7\lab7-SCHEMATIC1-Sim.sim ] 

** Creating circuit file "lab7-SCHEMATIC1-Sim.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 25ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\lab7-SCHEMATIC1.net" 


.END
