** Profile: "SCHEMATIC1-as"  [ F:\NUST\Semester 1\Linear Circuit Analysis\Labs\PSpice\short-SCHEMATIC1-as.sim ] 

** Creating circuit file "short-SCHEMATIC1-as.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\short-SCHEMATIC1.net" 


.END
